library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package cartram_comp is
	component cartram
	Port (
		RST : in STD_LOGIC;
		CLK : in  STD_LOGIC;
		ADDR : in STD_LOGIC_VECTOR(15 downto 0);
		RD_D : out STD_LOGIC_VECTOR(7 downto 0);
		WR_D : in STD_LOGIC_VECTOR(7 downto 0);
		OE : in STD_LOGIC;
		WR : in STD_LOGIC);
	end component;
end package;


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

library UNISIM;
use UNISIM.VComponents.all;

use work.types_comp.all;

entity cartram is
	Port (
		RST : in STD_LOGIC;
		CLK : in  STD_LOGIC;
		ADDR : in STD_LOGIC_VECTOR(15 downto 0);
		RD_D : out STD_LOGIC_VECTOR(7 downto 0);
		WR_D : in STD_LOGIC_VECTOR(7 downto 0);
		OE : in STD_LOGIC;
		WR : in STD_LOGIC);
end cartram;

architecture DataPath of cartram is

	signal in00, in08, in09 : ram_in;
	signal out00, out08, out09 : ram_out;

begin

	in00.addr <= ADDR(10 downto 0) & "000";
	in00.idata <= (others => '0');
	in00.ipar <= (others => '0');
	in00.wen <= (others => '0');  -- program ROM

	in08.addr <= ADDR(10 downto 0) & "000";
	in08.idata <= (others => '0');
	in08.ipar <= (others => '0');
	in08.wen <= (others => '0');  -- program ROM

	in09.addr <= ADDR(10 downto 0) & "000";
	in09.idata <= (others => '0');
	in09.ipar <= (others => '0');
	in09.wen <= (others => '0');  -- program ROM

	RD_D <= "ZZZZZZZZ"              WHEN OE = '0' ELSE
			out00.odata(7 downto 0) WHEN ADDR(15 downto 11) = "00000" ELSE  -- 0000-07FF
			out08.odata(7 downto 0) WHEN ADDR(15 downto 11) = "01000" ELSE  -- 4000-47FF
			out09.odata(7 downto 0) WHEN ADDR(15 downto 11) = "01001" ELSE  -- 4800-4FFF
	        "ZZZZZZZZ";

	ram00 : RAMB16BWER
	generic map (
		SIM_DEVICE => "SPARTAN6",
		DATA_WIDTH_A => 9,
		DATA_WIDTH_B => 9,
		WRITE_MODE_A => "WRITE_FIRST",
		WRITE_MODE_B => "WRITE_FIRST",
INIT_00 => X"0000000000c42cc30000000000c42cc30000000000c42cc30000000000c42cc3",
INIT_01 => X"0000000000c42cc30000000000c42cc30000000000c42cc30000000000c42cc3",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"e66eccdc0e0089881f1108000d000c00830073030b000dcc6666edce0213c300",
INIT_09 => X"474e494d49545f5254534e493e33b9bb9f99dcddccec0e6e6367bbbb99d9dddd",
INIT_0a => X"0000000000000000000000000000000050e7af00000000000100000080000000",
INIT_0b => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0c => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0d => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0e => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0f => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"000000000000000200c3400021c000c378f7200d14fb201c122a100ec0001147",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1a => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1b => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1c => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1d => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1e => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1f => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2a => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2b => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2c => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2d => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2e => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2f => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3a => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3b => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3c => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3d => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3e => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3f => X"0000000000000000000000000000000000000000000000000000000000000000",
		-- DOA_REG/DOB_REG: Optional output register (0 or 1)
		DOA_REG => 0,
		DOB_REG => 0,
		-- EN_RSTRAM_A/EN_RSTRAM_B: Enable/disable RST
		EN_RSTRAM_A => TRUE,
		EN_RSTRAM_B => TRUE,
		-- INIT_A/INIT_B: Initial values on output port
		INIT_A => X"000000000",
		INIT_B => X"000000000",
		-- RSTTYPE: "SYNC" or "ASYNC"
		RSTTYPE => "SYNC",
		-- RST_PRIORITY_A/RST_PRIORITY_B: "CE" or "SR"
		RST_PRIORITY_A => "CE",
		RST_PRIORITY_B => "CE",
		-- SIM_COLLISION_CHECK: Collision check enable "ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE"
		SIM_COLLISION_CHECK => "ALL",
		-- SIM_DEVICE: Must be set to "SPARTAN6" for proper simulation behavior
		-- SRVAL_A/SRVAL_B: Set/Reset value for RAM output
		SRVAL_A => X"000000000",
		SRVAL_B => X"000000000"
	)
	port map (
		-- Port A
		DOA => out00.odata,
		DOPA => out00.opar,
		ADDRA => in00.addr,
		CLKA => CLK,
		ENA => '1',
		REGCEA => '0',
		RSTA => RST,
		WEA => in00.wen,
		DIA => in00.idata,
		DIPA => in00.ipar,
		-- Port B
		ADDRB => "00" & X"000",   -- 14-bit input: B port address input
		CLKB => '0',	  -- 1-bit input: B port clock input
		ENB => '0',	   -- 1-bit input: B port enable input
		REGCEB => '0',	-- 1-bit input: B port register clock enable input
		RSTB => '0',	  -- 1-bit input: B port register set/reset input
		WEB => "0000",	-- 4-bit input: Port B byte-wide write enable input
		DIB => X"00000000",	   -- 32-bit input: B port data input
		DIPB => "0000"	-- 4-bit input: B port parity input
	);

	ram08 : RAMB16BWER
	generic map (
		SIM_DEVICE => "SPARTAN6",
		DATA_WIDTH_A => 9,
		DATA_WIDTH_B => 9,
		WRITE_MODE_A => "WRITE_FIRST",
		WRITE_MODE_B => "WRITE_FIRST",
INIT_00 => X"f5c8b7c9f6203df1c003cddf3ef5c8b7c900c8d001ce00301ffc3005d6c220c3",
INIT_01 => X"000000000000c9f1c003cd7dc010cd7cf5c9f1203df1c003cdd43ec012cdff3e",
INIT_02 => X"8321e5d5c5f5c983e082e081e080e0ff3e0018c9000000000000000000000000",
INIT_03 => X"5783ee7a4fb8ee7947edee785f10301f1acb19cb38cb0826ae2d562d4e2d46ff",
INIT_04 => X"18c93e0418d803ea7cd802ea7dc9f1c1d1e1702c712c7222ff26e4202520ee7b",
INIT_05 => X"d801cd0a3ef5c9f1d801cd203ef5c9f1d801cdc05ac40afef5c9d801eac33e02",
INIT_06 => X"cdc123cdc11dcdc113cdc0eecdc9f1f920b72ac0a7cd0318f5e9c0c7cde1c9f1",
INIT_07 => X"f5e51878f5c9c1c0ffcdc1f5c5f1c129cdf5c9f1d801cd203ec129cdf5c9c0ba",
INIT_08 => X"42c5f5c718c179c129cd78c5f5d1187df5d5187cf5d9187bf5dd187af5e11879",
INIT_09 => X"d801c330c607c602380afe0fe6f1c133cd37cbf5c05acdec184d44c5f5f2184b",
INIT_0a => X"042f06c9f1c1c0a7cd30c6c15dcd0a0ec15dd4b9640e0b380afec5f50c18c5f5",
INIT_0b => X"cde5c9f1d806ea7cd805ea7dd804ea2a2323f5e5e1c979c0a7cd784f81fc3091",
INIT_0c => X"fac26bc3003ee100646573736150c0c2cde5c0bacdc9c04dcde100ff0218c16b",
INIT_0d => X"d806fa6fd805fac26bc3003ee100656e6f44c0c2cde50f18e3283d05283cd804",
INIT_0e => X"2f81f0f52f80f0f5c26bc300ce01fed804fac0bacdc0c7cdc0bacd0928b77e67",
INIT_0f => X"81f01220bb80f0c9f1c0e3cdf1c129cdf1c129cdf1c129cd2f83f0f52f82f0f5",
INIT_10 => X"c9f720b1780bc05acd2ac1b9c3c1d8cdc04fc30320b883f00820b982f00d20ba",
INIT_11 => X"3e25e0ff3e26e0803e26e0003effe0003e0fe0003e07e0003ed800eadfff31f3",
INIT_12 => X"cdcd3ec012cdff3ec01fcd033ef5c04fcdc877cdc17ecdc093cdc88f2124e077",
INIT_13 => X"01fef1c0a1cdc0bacdf5c8a6c3f1c276cdf5dfff31c26bc3003ec300cdf1c003",
INIT_14 => X"cde100232064656c696146c0c2cde5c9e1000a64656c696146c0c2cde50e20d8",
INIT_15 => X"3ef505e0ec3e0fe0003e07e0053e06e0003effe004e6fff0f3f5c9c0bacdc144",
INIT_16 => X"c9f1f820b705f005e0aff5c9f1c1b9ca04e60ff0c1b9c204e60ff0f1c003cd29",
INIT_17 => X"c9f720b71b05f005e0af5f12cb8712cb8705d605f00016c9d10ad67bc2e9cdd5",
INIT_18 => X"c8b7c2e0cdc2d5cdc19fc3c3a3cdc348cde100000218c16bcde5c318cdc2a6cd",
INIT_19 => X"65706f7270206b726f77202074276e73656f642072656d6954021e18c16bcde5",
INIT_1a => X"e6d800fa0620c7e62f7dc9f5202cc356c400fe7eca26002ec1b9c3e100796c72",
INIT_1b => X"c8bac8becb26c384cd5f2f7bc3decd570428be0016c384cd5ff8c608e67dc004",
INIT_1c => X"c404cd7b22d83e22263e05280d003e0b280d22d820217d4ec926e5d5c9c3decd",
INIT_1d => X"0120bec3cecdff1e0920bec3cecd001ec9f7202cc3b0c400fe7ecc0021c9d1e1",
INIT_1e => X"7df5c9e1c404cdd820eacb3e22d821217de5c9c3decde100204243c0c2cde5c9",
INIT_1f => X"0218c16bcde5c0a7cd203ec144cd7ec0a7cd2d3ec144cdf1c0a7cd3a3ec129cd",
INIT_20 => X"2611d82601c5d81e0877d828eac43e22d827ea2c3ed826ea22c33e4fc9e10001",
INIT_21 => X"28b17803fb1e01c5c918d6c2e0cdf9e1d81e31f3d820c3e5f1c2d5cdd82621d8",
INIT_22 => X"c4cd000e820021c47dcd203ec48bc410e6d800fac4eccdc9c1f52090fe44f006",
INIT_23 => X"9800215c18c532cdd81deaf83ed81cea003ed81bea143ec4c4cdff0e8a0021c4",
INIT_24 => X"e0003e69e0003e69e07f3e69e0ff3e100668e0803ec9f8200524fc202c770406",
INIT_25 => X"003ec47dcd003eff4fea013edd200569e0003e69e0003e69e0003e69e0003e69",
INIT_26 => X"e0913ec438cdf5c9f12005c1f820052222a9131a0806c56006c57711c9ff4fea",
INIT_27 => X"d81cea80e6803e0218afc9f140e0113ec438cdf5c556c347e0e43e43e0003e40",
INIT_28 => X"e1776e352db6f1f5c522cd0a2820fef1092007fe2ad81b21f5e51d280afef5c9",
INIT_29 => X"1a21203ed81dea08c6d81dfae5c5c556c3c55fcdc532cdc55fcdc438cdf5c9f1",
INIT_2a => X"d5c9f142e088d6d81dfac55fcdc438cdf5c9c1e1d81bea1b3efc2005321406d8",
INIT_2b => X"180000000000000000c9d1e1f82007fe7b221a1dd81b11292926266fd81dfae5",
INIT_2c => X"6600187c063c603e1800006cfe6c6cfe6c00000000006c6c6c00180018181818",
INIT_2d => X"70000e1c1818181c0e00000000000c0c0c003b666f381c361c0086c66030186c",
INIT_2e => X"006030300000000000000018187e1818000000663cff3c660000703818181838",
INIT_2f => X"18003c6666766e663c00406030180c06020060600000000000000000007e0000",
INIT_30 => X"7e000c0c7e6c3c1c0c003c66060c180c7e007e30180c06663c007e1818181838",
INIT_31 => X"3c003c66663c66663c00303030180c067e003c66667c60603c003c6606067c60",
INIT_32 => X"00000c18306030180c0030181800181800000018180018180000380c063e6666",
INIT_33 => X"18003e606e6a6e663c001800180c06663c0030180c060c183000007e00007e00",
INIT_34 => X"7e00786c6666666c78003c66606060663c007c66667c66667c0066667e66663c",
INIT_35 => X"3c006666667e666666003e66666e60603e006060607c60607e007e60607c6060",
INIT_36 => X"c6007e60606060606000666c7870786c66003c660606060606003c1818181818",
INIT_37 => X"3c006060607c66667c003c66666666663c0066666e7e7e766600c6c6c6d6feee",
INIT_38 => X"66001818181818187e003c66063c60663c0066666c7c66667c00366c76666666",
INIT_39 => X"660066663c183c666600c6eefed6c6c6c600183c3c66666666003e6666666666",
INIT_3a => X"780002060c18306040001e18181818181e007e6030180c067e001818183c6666",
INIT_3b => X"0000000000003060c0fe0000000000000000000000c66c381000781818181818",
INIT_3c => X"00003e6666663e0606003c6060603c0000007c6666667c6060003e663e063c00",
INIT_3d => X"1800666666667c60607c063e66663e000000303030307c301c003c607e663c00",
INIT_3e => X"00003c18181818183800666c786c6660607018181818180018003c1818183800",
INIT_3f => X"00607c6666667c0000003c6666663c000000666666667c000000c6c6d6feec00",
		-- DOA_REG/DOB_REG: Optional output register (0 or 1)
		DOA_REG => 0,
		DOB_REG => 0,
		-- EN_RSTRAM_A/EN_RSTRAM_B: Enable/disable RST
		EN_RSTRAM_A => TRUE,
		EN_RSTRAM_B => TRUE,
		-- INIT_A/INIT_B: Initial values on output port
		INIT_A => X"000000000",
		INIT_B => X"000000000",
		-- RSTTYPE: "SYNC" or "ASYNC"
		RSTTYPE => "SYNC",
		-- RST_PRIORITY_A/RST_PRIORITY_B: "CE" or "SR"
		RST_PRIORITY_A => "CE",
		RST_PRIORITY_B => "CE",
		-- SIM_COLLISION_CHECK: Collision check enable "ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE"
		SIM_COLLISION_CHECK => "ALL",
		-- SIM_DEVICE: Must be set to "SPARTAN6" for proper simulation behavior
		-- SRVAL_A/SRVAL_B: Set/Reset value for RAM output
		SRVAL_A => X"000000000",
		SRVAL_B => X"000000000"
	)
	port map (
		-- Port A
		DOA => out08.odata,
		DOPA => out08.opar,
		ADDRA => in08.addr,
		CLKA => CLK,
		ENA => '1',
		REGCEA => '0',
		RSTA => RST,
		WEA => in08.wen,
		DIA => in08.idata,
		DIPA => in08.ipar,
		-- Port B
		ADDRB => "00" & X"000",   -- 14-bit input: B port address input
		CLKB => '0',	  -- 1-bit input: B port clock input
		ENB => '0',	   -- 1-bit input: B port enable input
		REGCEB => '0',	-- 1-bit input: B port register clock enable input
		RSTB => '0',	  -- 1-bit input: B port register set/reset input
		WEB => "0000",	-- 4-bit input: Port B byte-wide write enable input
		DIB => X"00000000",	   -- 32-bit input: B port data input
		DIPB => "0000"	-- 4-bit input: B port parity input
	);

	ram09 : RAMB16BWER
	generic map (
		SIM_DEVICE => "SPARTAN6",
		DATA_WIDTH_A => 9,
		DATA_WIDTH_B => 9,
		WRITE_MODE_A => "WRITE_FIRST",
		WRITE_MODE_B => "WRITE_FIRST",
INIT_00 => X"00000e1818187e1800007c063c603e000000606060667c0000063e6666663e00",
INIT_01 => X"0000663c183c660000006c7cd6c6c6000000183c6666660000003e6666666600",
INIT_02 => X"700018181818181818000e18183018180e007e30180c7e00007c063e66666600",
INIT_03 => X"6e69c0c2cde5c449cd000000000000000000000c9ef2600000007018180c1818",
INIT_04 => X"03cdd83ec012cd083ef502e0813e01e0f5c9e1000a0a676e696d69745f727473",
INIT_05 => X"00000000000000000000000000c9fe1826e0003ec8b2cdc4d9cdc501c3f1f1c0",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0102010101010102010201010101030001020101010101030102010101010301",
INIT_09 => X"0102010101010102010201010101030201020101010101020102010101010302",
INIT_0a => X"0101010101010101010101010101010101010101010101010101010101010101",
INIT_0b => X"0101010101010101010101010101010101010101010101010101010101010101",
INIT_0c => X"0101010101010101010101010101010101010101010101010101010101010101",
INIT_0d => X"0101010101010101010101010101010101010101010101010101010101010101",
INIT_0e => X"0102000300030101010201030003010101020303000301010102010303030101",
INIT_0f => X"0102000001030102010201000101010201020000000301020102010000010102",
INIT_10 => X"0102010102020203010201010202030001020101020202050102010102020301",
INIT_11 => X"0102010102020202010303030202030201020101020202020102010102020302",
INIT_12 => X"0102010101010101010201010101010101020101010101010102010101010101",
INIT_13 => X"0102010101010101020002020202020201020101010101010102010101010101",
INIT_14 => X"0102010101010101010201010101010101020101010101010102010101010101",
INIT_15 => X"0102010101010101010201010101010101020101010101010102010101010101",
INIT_16 => X"0402000300030402040204030003030204020603000304020402040304030302",
INIT_17 => X"0402000001040203040204000102030304020000000401040402040000020303",
INIT_18 => X"0102010102020203010201010202030001020101020202050102010102020301",
INIT_19 => X"0102010102020203010303030202030301020101020202030102010102020303",
INIT_1a => X"0102010101010101010201010101010101020101010101010102010101010101",
INIT_1b => X"0102010101010101020002020202020201020101010101010102010101010101",
INIT_1c => X"0102010101010101010201010101010101020101010101010102010101010101",
INIT_1d => X"0102010101010101010201010101010101020101010101010102010101010101",
INIT_1e => X"0402000600040405040204060004030504020606000404050402040604040305",
INIT_1f => X"0402000001040203040204000102030304020000000401040402040000020303",
INIT_20 => X"0204020202020202020402020202020202040202020202020204020202020202",
INIT_21 => X"0204020202020202020402020202020202040202020202020204020202020202",
INIT_22 => X"0203020202020202020302020202020202030202020202020203020202020202",
INIT_23 => X"0203020202020202020302020202020202030202020202020203020202020202",
INIT_24 => X"0204020202020202020402020202020202040202020202020204020202020202",
INIT_25 => X"0204020202020202020402020202020202040202020202020204020202020202",
INIT_26 => X"0204020202020202020402020202020202040202020202020204020202020202",
INIT_27 => X"0204020202020202020402020202020202040202020202020204020202020202",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2a => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2b => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2c => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2d => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2e => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2f => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3a => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3b => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3c => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3d => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3e => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3f => X"0000000000000000000000000000000000000000000000000000000000000000",
		-- DOA_REG/DOB_REG: Optional output register (0 or 1)
		DOA_REG => 0,
		DOB_REG => 0,
		-- EN_RSTRAM_A/EN_RSTRAM_B: Enable/disable RST
		EN_RSTRAM_A => TRUE,
		EN_RSTRAM_B => TRUE,
		-- INIT_A/INIT_B: Initial values on output port
		INIT_A => X"000000000",
		INIT_B => X"000000000",
		-- RSTTYPE: "SYNC" or "ASYNC"
		RSTTYPE => "SYNC",
		-- RST_PRIORITY_A/RST_PRIORITY_B: "CE" or "SR"
		RST_PRIORITY_A => "CE",
		RST_PRIORITY_B => "CE",
		-- SIM_COLLISION_CHECK: Collision check enable "ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE"
		SIM_COLLISION_CHECK => "ALL",
		-- SIM_DEVICE: Must be set to "SPARTAN6" for proper simulation behavior
		-- SRVAL_A/SRVAL_B: Set/Reset value for RAM output
		SRVAL_A => X"000000000",
		SRVAL_B => X"000000000"
	)
	port map (
		-- Port A
		DOA => out09.odata,
		DOPA => out09.opar,
		ADDRA => in09.addr,
		CLKA => CLK,
		ENA => '1',
		REGCEA => '0',
		RSTA => RST,
		WEA => in09.wen,
		DIA => in09.idata,
		DIPA => in09.ipar,
		-- Port B
		ADDRB => "00" & X"000",   -- 14-bit input: B port address input
		CLKB => '0',	  -- 1-bit input: B port clock input
		ENB => '0',	   -- 1-bit input: B port enable input
		REGCEB => '0',	-- 1-bit input: B port register clock enable input
		RSTB => '0',	  -- 1-bit input: B port register set/reset input
		WEB => "0000",	-- 4-bit input: Port B byte-wide write enable input
		DIB => X"00000000",	   -- 32-bit input: B port data input
		DIPB => "0000"	-- 4-bit input: B port parity input
	);

end DataPath;
